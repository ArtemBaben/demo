`timescale 1ns / 1ps
`default_nettype none
/*
//////////////////////////////////////////////////////////////////////////////////
// Company 		:  	RNIIRS
// Engineer		:  	Babenko Artem
// 
// Description  :	binary_offset2Twos_complement module 
//
//
//
//
/////////////////////////////////////////////////////////////////////////////////
*/
module bo2tc
#(
parameter 			PORTS								= 8				
)
(
// system_interface
input	wire		[(PORTS-1):0][7:0]					DATA_IN		,
output	wire		[(PORTS-1):0][7:0]					DATA_OUT	
);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Wires and regs
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
genvar 			i;

generate
for (i=0;i<PORTS;i=i+1) begin : binary_offset2twos_complement
	assign DATA_OUT[i] = {~DATA_IN[i][7],DATA_IN[i][6:0]};
end
endgenerate




endmodule
`default_nettype wire